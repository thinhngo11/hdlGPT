module evenodd (output Y, input A, B, B, C);
  assign Y = A ^ B ^ C ^ D;
endmodule
