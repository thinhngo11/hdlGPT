interface magnitude_comparator_if(input logic clk);
    logic [3:0] A;
    logic [3:0] B;
    logic A_greater;
    logic A_equal;
    logic A_less;
endinterface
